module structural (
    input wire A,
    input wire B,
    output wire C
);
and and_test(C, A, B);
endmodule